`timescale 1ns / 1ps
`default_nettype none

module jojo(
  output logic [159:0][5:0] jonathan
);
  assign jonathan[0] = 6'b0_00000;
  assign jonathan[1] = 6'b0_00000;
  assign jonathan[2] = 6'b0_00000;
  assign jonathan[3] = 6'b0_00000;
  assign jonathan[4] = 6'b0_00000;
  assign jonathan[5] = 6'b0_00000;
  assign jonathan[6] = 6'b1_00010;
  assign jonathan[7] = 6'b1_00101;

  assign jonathan[8] = 6'b1_01001;
  assign jonathan[9] = 6'b1_01001;
  assign jonathan[10] = 6'b1_01110;
  assign jonathan[11] = 6'b1_01110;
  assign jonathan[12] = 6'b1_01100;
  assign jonathan[13] = 6'b1_01100;
  assign jonathan[14] = 6'b1_00111;
  assign jonathan[15] = 6'b1_00111;
  
  assign jonathan[16] = 6'b1_00101;
  assign jonathan[17] = 6'b1_00111;
  assign jonathan[18] = 6'b1_01001;
  assign jonathan[19] = 6'b1_01001;
  assign jonathan[20] = 6'b1_01001;
  assign jonathan[21] = 6'b1_01001;
  assign jonathan[22] = 6'b1_01001;
  assign jonathan[23] = 6'b1_00111;
  
  assign jonathan[24] = 6'b1_00101;
  assign jonathan[25] = 6'b1_00101;
  assign jonathan[26] = 6'b1_01001;
  assign jonathan[27] = 6'b1_01001;
  assign jonathan[28] = 6'b1_00111;
  assign jonathan[29] = 6'b1_00111;
  assign jonathan[30] = 6'b1_00100;
  assign jonathan[31] = 6'b1_00100;

  assign jonathan[32] = 6'b1_00010;
  assign jonathan[33] = 6'b1_00010;
  assign jonathan[34] = 6'b1_00010;
  assign jonathan[35] = 6'b1_00010;
  assign jonathan[36] = 6'b1_00010;
  assign jonathan[37] = 6'b1_00010;
  assign jonathan[38] = 6'b1_00010;
  assign jonathan[39] = 6'b1_00101;

  assign jonathan[40] = 6'b1_01001;
  assign jonathan[41] = 6'b1_01001;
  assign jonathan[42] = 6'b1_01110;
  assign jonathan[43] = 6'b1_01110;
  assign jonathan[44] = 6'b1_01100;
  assign jonathan[45] = 6'b1_01100;
  assign jonathan[46] = 6'b1_00111;
  assign jonathan[47] = 6'b1_00111;

  assign jonathan[48] = 6'b1_10000;
  assign jonathan[49] = 6'b1_10000;
  assign jonathan[50] = 6'b1_10001;
  assign jonathan[51] = 6'b1_10000;
  assign jonathan[52] = 6'b1_01110;
  assign jonathan[53] = 6'b1_01110;
  assign jonathan[54] = 6'b1_01100;
  assign jonathan[55] = 6'b1_01010;

  assign jonathan[56] = 6'b1_01001;
  assign jonathan[57] = 6'b1_01001;
  assign jonathan[58] = 6'b1_00111;
  assign jonathan[59] = 6'b1_00101;
  assign jonathan[60] = 6'b1_00111;
  assign jonathan[61] = 6'b1_00111;
  assign jonathan[62] = 6'b1_00100;
  assign jonathan[63] = 6'b1_00100;

  assign jonathan[64] = 6'b1_00010;
  assign jonathan[65] = 6'b1_00010;
  assign jonathan[66] = 6'b1_00010;
  assign jonathan[67] = 6'b1_00010;
  assign jonathan[68] = 6'b1_00010;
  assign jonathan[69] = 6'b1_00010;//'NICE!' - Joseph jonathan
  assign jonathan[70] = 6'b1_00010;
  assign jonathan[71] = 6'b1_00010;
  assign jonathan[159:72] = 0;
endmodule


`default_nettype wire

